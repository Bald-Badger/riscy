`include "../../opcode.vh"

module pc_adder_tb (

);
	
endmodule
