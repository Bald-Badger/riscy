import defines::*;
import mem_defines::*;

module cache(
	input logic		clk,
	input logic		rst_n,
	input tag_t		tag,
	input offset_t	offset,
	input data_t	data_in,
);
	
endmodule : cache
