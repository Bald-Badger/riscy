// functional model of a sram inetrface

module sram(
	
);
	
endmodule : sram
