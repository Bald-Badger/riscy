bind memory memory_sva check_memory(
    clk,
	clk_100m,
	clk_100m_shift,
	rst_n,
	addr,
	data_in_raw,
	mem_mem_fwd_data,
	fwd_m2m,
	instr,
	data_out,
	sdram_init_done,
	done,
	sdram_clk, 
	sdram_cke,
	sdram_cs_n,   
	sdram_ras_n,
	sdram_cas_n,
	sdram_we_n,
	sdram_ba,
	sdram_addr,
	sdram_data,
	sdram_dqm
);