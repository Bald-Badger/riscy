`include "../../opcode.vh"

module extend (
    
);
    
endmodule