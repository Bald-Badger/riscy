module pref (
	
);
	
endmodule : pref
