`include "../opcode.svh"
`include "./alu_define.svh"

module alu_tb ();

instr_t instr;
data_t a_in, b_in, c_out;



endmodule
