package pref_defines;
import defines::*;
import mem_defines::*;

`ifndef _pref_defines_
`define _pref_defines_


// defined in mem_defines
// localparam	MAX_PHY_MEM			= 32'h01ff_ffff
// localparam	MMIO_BASE			= 32'h0200_0000

`endif
endpackage : pref_defines
