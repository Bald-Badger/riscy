import defines::*;

module hazzard_ctrl (
	// input signal
	input instr_t instr_f,
	input instr_t instr_d,
	input instr_t instr_x,
	input instr_t instr_m,
	input instr_t instr_w,

	input logic ex_mem_wr_rd,
	input logic mem_wb_wr_rd,

	input branch_take_t branch_predict,
	input branch_take_t branch_actual,

	// forwarding signal
	output fwd_sel_t fwd_a,
	output fwd_sel_t fwd_b,
	output fwd_sel_t fwd_m2m,

	output branch_fwd_t fwd_rs1,
	output branch_fwd_t fwd_rs2,

	// stall signal
	output logic stall_if_id,
	output logic stall_id_ex,
	output logic stall_ex_mem,
	output logic stall_mem_wb,

	// flush signal
	output logic flush_if_id,
	output logic flush_id_ex,
	output logic flush_ex_mem,
	output logic flush_mem_wb
);
	

	r_t id_ex_rs1, id_ex_rs2, ex_mem_rs2, ex_mem_rd, mem_wb_rd;
	logic mem_store;
	always_comb begin : input_sig
		id_ex_rs1 = instr_x.rs1;
		id_ex_rs2 = instr_x.rs2;
		ex_mem_rs2 = instr_m.rs2;
		ex_mem_rd = instr_m.rd;
		mem_wb_rd = instr_w.rd;
		mem_store = (instr_m.opcode == STORE);
	end


	logic hazzard_1a, hazzard_1b, hazzard_2a, hazzard_2b, hazzard_3;

	always_comb begin : data_hazzard_detect

		hazzard_1a =	(ex_mem_wr_rd) &&
						(ex_mem_rd != X0) &&
						(ex_mem_rd == id_ex_rs1);
	
		hazzard_1b =	(ex_mem_wr_rd) &&
						(ex_mem_rd != X0) &&
						(ex_mem_rd == id_ex_rs2);

		hazzard_2a =	(mem_wb_wr_rd) &&
						(mem_wb_rd != X0) &&
						(!(ex_mem_wr_rd && 
							(ex_mem_wr_rd != X0) &&
							(ex_mem_wr_rd == id_ex_rs1))) &&
						(mem_wb_rd == id_ex_rs1);
		
		hazzard_2b =	(mem_wb_wr_rd) &&
						(mem_wb_rd != X0) &&
						(!(ex_mem_wr_rd && 
							(ex_mem_wr_rd != X0) &&
							(ex_mem_wr_rd == id_ex_rs1))) &&
						(mem_wb_rd == id_ex_rs2);
	
		hazzard_3 =		(mem_store) &&
						(ex_mem_rd != X0) && 
						(mem_wb_rd == ex_mem_rs2);

	end


	always_comb begin : forward_sig_assign

		fwd_a =	hazzard_1a ? EX_EX_FWD_SEL :
				hazzard_2a ? MEM_EX_FWD_SEL :
				RS_SEL;

		fwd_b = hazzard_1b ? EX_EX_FWD_SEL :
				hazzard_2b ? MEM_EX_FWD_SEL :
				RS_SEL;
		
		fwd_m2m = hazzard_3 ? MEM_MEM_FWD_SEL : RS_SEL;

	end

	always_comb begin : control_hazzard_detect
		
	end

	
	
endmodule : hazzard_ctrl
