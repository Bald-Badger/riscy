`include "../opcode.svh"

module alu (
	
);
	
endmodule
