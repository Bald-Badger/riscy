import defines::*;

module pref ();
	
endmodule : pref
