import defines::*;
import mem_defines::*;

module mem_ctrl (
	
);
	
endmodule: mem_ctrl
