`include "../opcode.svh"

module ex_mux (
	
);
	
endmodule
