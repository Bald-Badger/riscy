`include "./opcode.svh"
`timescale 1ns/1ns

module proc_hier_tb ();
	
	proc_hier proc_hier_inst();

endmodule
